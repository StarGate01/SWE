(
        netcdf foo { // example netCDF specification in CDL
        dimensions:
            lat = 10, lon = 5, time = unlimited;
        variables:
            int lat(lat), lon(lon), time(time);
            float z(time,lat,lon), t(lat,lon);
            lat:units = "degrees_north";
            lon:units = "degrees_east";
            time:units = "seconds";
            z:valid_range = 0., 5000.;
            :test = "global value";
        data:
       lat = 0, 10, 20, 30, 40, 50, 60, 70, 80, 90;
    invalid data
)